//Universidad del Valle de Guatemala
//Gerardo Fuentes
// 19389

module testbench();

  reg t1, t2, t3;
  wire s1, s2, s3, s4, s5, s6;

  
